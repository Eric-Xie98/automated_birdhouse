module and_32bit(o, A, B);

    input [31:0] A, B;
    output [31:0] o;

    and a0(o[0], A[0], B[0]);
    and a1(o[1], A[1], B[1]);
    and a2(o[2], A[2], B[2]);
    and a3(o[3], A[3], B[3]);
    and a4(o[4], A[4], B[4]);
    and a5(o[5], A[5], B[5]);
    and a6(o[6], A[6], B[6]);
    and a7(o[7], A[7], B[7]);
    and a8(o[8], A[8], B[8]);
    and a9(o[9], A[9], B[9]);
    and a10(o[10], A[10], B[10]);
    and a11(o[11], A[11], B[11]);
    and a12(o[12], A[12], B[12]);
    and a13(o[13], A[13], B[13]);
    and a14(o[14], A[14], B[14]);
    and a15(o[15], A[15], B[15]);
    and a16(o[16], A[16], B[16]);
    and a17(o[17], A[17], B[17]);
    and a18(o[18], A[18], B[18]);
    and a19(o[19], A[19], B[19]);
    and a20(o[20], A[20], B[20]);
    and a21(o[21], A[21], B[21]);
    and a22(o[22], A[22], B[22]);
    and a23(o[23], A[23], B[23]);
    and a24(o[24], A[24], B[24]);
    and a25(o[25], A[25], B[25]);
    and a26(o[26], A[26], B[26]);
    and a27(o[27], A[27], B[27]);
    and a28(o[28], A[28], B[28]);
    and a29(o[29], A[29], B[29]);
    and a30(o[30], A[30], B[30]);
    and a31(o[31], A[31], B[31]);

endmodule